library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity WS2812B_driver is
	generic (
		max_pos : integer := 16
	);
	
	port (
		clk : in std_logic;
		enable : in std_logic;
		leds_line : out std_logic := '0';
		
		seq_sequence : out std_logic := '0';
		
		update_frame : in std_logic;
		
		program_led_number : buffer integer range 0 to max_pos-1;
		program_red_intensity : in integer range 0 to 255;
		program_blue_intensity : in integer range 0 to 255;
		program_green_intensity : in integer range 0 to 255
	);
end entity;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity NRZ_sequence is
	generic (
		duration_clk_counts : integer;
		code_0_high_duration_clk_counts : integer;
		code_1_high_duration_clk_counts : integer
	);
	
	port (
		clk : in std_logic;
		trigger : in std_logic;
		finished : in std_logic;
		bit_to_code : in std_logic;
		sequence : out std_logic := '0'
	);

end entity;

architecture behavior of NRZ_sequence is
	signal step : integer range 0 to duration_clk_counts := 0;
	signal is_start : std_logic := '0';
	
	signal stim_start : std_logic;
begin

	process(stim_start)
	begin
		if rising_edge(stim_start) then
			if trigger = '1' then
				is_start <= '1';
			else
				is_start <= '0';
			end if;
		end if;
	end process;

	process(clk)
	begin
		if rising_edge(clk) then
			if is_start = '1' then
			
				if step = duration_clk_counts then
					step <= 0;
				else
					step <= step + 1;
				end if;
			end if;
		end if;
	end process;
	
	stim_start <= '1' when (is_start = '0' and trigger = '1') or (trigger = '0' and is_start = '1' and step = 0) else '0';

	sequence <= '1' when ((bit_to_code = '0' and step <= 19) or (bit_to_code = '1' and step <= 39)) and is_start = '1' else '0';
	
end architecture;


architecture beh of WS2812B_driver is
	constant step_max : integer := 62;
	constant bit_proceed_max : integer := 23;

	signal step : integer range 0 to step_max;
	signal bit_proceed : integer range 0 to bit_proceed_max;

	constant WaitStart : std_logic_vector(0 to 1) := "00";
	constant SendLEDsData : std_logic_vector(0 to 1) := "01";
	constant ValidateSeq : std_logic_vector(0 to 1) := "10";
	
	signal stage : std_logic_vector(0 to 1) := WaitStart;
	
	signal seq_trigger : std_logic;
	signal seq_finished : std_logic;
	signal seq_bit_to_code : std_logic;
	
	constant HIGH_DURATION_FOR_CODE_1 : integer := 39;
	constant HIGH_DURATION_FOR_CODE_0 : integer := 19;
	
	function serial_state_led_line_for_color (
		step : integer range 0 to step_max;
		bit_proceed : integer range 0 to bit_proceed_max;
		
		green: integer range 0 to 255;
		red: integer range 0 to 255;
		blue: integer range 0 to 255
	) return std_logic is
		variable data :  std_logic_vector(0 to bit_proceed_max);
	begin
		data := std_logic_vector( to_unsigned( green, 8)) & std_logic_vector( to_unsigned( red, 8)) & std_logic_vector( to_unsigned( blue, 8));
	
		if data(bit_proceed) = '0' and step <= HIGH_DURATION_FOR_CODE_0 then
			return '1';
		elsif data(bit_proceed) = '1' and step <= HIGH_DURATION_FOR_CODE_1 then
			return '1';
		else
			return '0';
		end if;
	end function;
begin
	NRZ_sequence : entity work.NRZ_sequence
		generic map(
			duration_clk_counts => 62,
			code_1_high_duration_clk_counts => 39,
			code_0_high_duration_clk_counts => 19
		)
		port map (
			clk => clk,
			trigger => seq_trigger,
			finished => seq_finished,
			bit_to_code => seq_bit_to_code,
			sequence => leds_line
		);

	process(clk)
		variable data :  std_logic_vector(0 to bit_proceed_max);
	begin
	
		data := std_logic_vector( to_unsigned( program_green_intensity, 8)) & std_logic_vector( to_unsigned( program_red_intensity, 8)) & std_logic_vector( to_unsigned( program_blue_intensity, 8));
	
		if rising_edge(clk) then
			case stage is
				when WaitStart =>
					seq_trigger <= '0';
				
					if enable = '1' then
						seq_trigger <= '1';
						seq_bit_to_code <= data(bit_proceed);
						stage <= SendLEDsData;
					end if;		
				when SendLEDsData =>
					if step = step_max then
						step <= 0;
						
						if bit_proceed = bit_proceed_max then
							bit_proceed <= 0;
							seq_bit_to_code <= data(0);
							seq_trigger <= '1';
							
							if program_led_number = max_pos-1 then
								program_led_number <= 0;
								
								stage <= ValidateSeq;
							else
								program_led_number <= program_led_number + 1;
							end if;
						else
							seq_trigger <= '1';

							bit_proceed <= bit_proceed + 1;
							seq_bit_to_code <= data(bit_proceed + 1);
						end if;
					else
						step <= step + 1;
						
						seq_trigger <= '0';
					end if;
				
				when ValidateSeq =>
					if update_frame = '1' then
						seq_trigger <= '1';

						stage <= SendLEDsData;
					else
						seq_trigger <= '0';
					end if;

				when others =>
					--nothing todo
			end case;
		end if;

	end process;

end architecture;